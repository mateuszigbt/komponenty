   �     7   :  P     7   _registeredBookmarks  :  {"api/WyświetlanieDanych.Form1.html":["wrapper","autocollapse","logo","navbar","search","search-query","breadcrumb","sidetoggle","sidetoc","_content","Wy_wietlanieDanych_Form1","Wy_wietlanieDanych_Form1_syntax","constructors","Wy_wietlanieDanych_Form1__ctor_","Wy_wietlanieDanych_Form1__ctor","Wy_wietlanieDanych_Form1__ctor_System_Runtime_Serialization_SerializationInfo_System_Runtime_Serialization_StreamingContext_","methods","Wy_wietlanieDanych_Form1_Dispose_","Wy_wietlanieDanych_Form1_Dispose_System_Boolean_","Wy_wietlanieDanych_Form1_GetObjectData_","Wy_wietlanieDanych_Form1_GetObjectData_System_Runtime_Serialization_SerializationInfo_System_Runtime_Serialization_StreamingContext_","implements","affix","viewport","title","generator"],"api/WyświetlanieDanych.Form2.html":["wrapper","autocollapse","logo","navbar","search","search-query","breadcrumb","sidetoggle","sidetoc","_content","Wy_wietlanieDanych_Form2","Wy_wietlanieDanych_Form2_syntax","constructors","Wy_wietlanieDanych_Form2__ctor_","Wy_wietlanieDanych_Form2__ctor","fields","Wy_wietlanieDanych_Form2_chart1","Wy_wietlanieDanych_Form2_circularProgressBar1","Wy_wietlanieDanych_Form2_trackBar1","properties","Wy_wietlanieDanych_Form2_Name1_","Wy_wietlanieDanych_Form2_Name1","Wy_wietlanieDanych_Form2_Name2_","Wy_wietlanieDanych_Form2_Name2","Wy_wietlanieDanych_Form2_Name3_","Wy_wietlanieDanych_Form2_Name3","methods","Wy_wietlanieDanych_Form2_Dispose_","Wy_wietlanieDanych_Form2_Dispose_System_Boolean_","implements","affix","viewport","title","generator"],"api/WyświetlanieDanych.KomponentOdbieranie.html":["wrapper","autocollapse","logo","navbar","search","search-query","breadcrumb","sidetoggle","sidetoc","_content","Wy_wietlanieDanych_KomponentOdbieranie","classes","affix","viewport","title","generator"],"api/WyświetlanieDanych.OdbieranieDanych.html":["wrapper","autocollapse","logo","navbar","search","search-query","breadcrumb","sidetoggle","sidetoc","_content","Wy_wietlanieDanych_OdbieranieDanych","Wy_wietlanieDanych_OdbieranieDanych_syntax","constructors","Wy_wietlanieDanych_OdbieranieDanych__ctor_","Wy_wietlanieDanych_OdbieranieDanych__ctor_System_String_","properties","Wy_wietlanieDanych_OdbieranieDanych_dateTime_","Wy_wietlanieDanych_OdbieranieDanych_dateTime","Wy_wietlanieDanych_OdbieranieDanych_PortName_","Wy_wietlanieDanych_OdbieranieDanych_PortName","Wy_wietlanieDanych_OdbieranieDanych_Wartosci_","Wy_wietlanieDanych_OdbieranieDanych_Wartosci","methods","Wy_wietlanieDanych_OdbieranieDanych_serialPort_DataRecived_","Wy_wietlanieDanych_OdbieranieDanych_serialPort_DataRecived_System_Object_System_IO_Ports_SerialDataReceivedEventArgs_","events","Wy_wietlanieDanych_OdbieranieDanych_DataReceived","affix","viewport","title","generator"],"api/WyświetlanieDanych.KomponentOdbieranie.Run_odbieranie.html":["wrapper","autocollapse","logo","navbar","search","search-query","breadcrumb","sidetoggle","sidetoc","_content","Wy_wietlanieDanych_KomponentOdbieranie_Run_odbieranie","Wy_wietlanieDanych_KomponentOdbieranie_Run_odbieranie_syntax","methods","Wy_wietlanieDanych_KomponentOdbieranie_Run_odbieranie_Main_","Wy_wietlanieDanych_KomponentOdbieranie_Run_odbieranie_Main","affix","viewport","title","generator"],"articles/intro.html":["wrapper","autocollapse","logo","navbar","search","search-query","breadcrumb","sidetoggle","sidetoc","_content","add-your-introductions-here","affix","viewport","title","generator"],"index.html":["wrapper","autocollapse","logo","navbar","search","search-query","breadcrumb","_content","this-is-the-homepage","quick-start-notes","affix","viewport","title","generator"],"api/index.html":["wrapper","autocollapse","logo","navbar","search","search-query","breadcrumb","sidetoggle","sidetoc","_content","placeholder","affix","viewport","title","generator"],"api/WyświetlanieDanych.html":["wrapper","autocollapse","logo","navbar","search","search-query","breadcrumb","sidetoggle","sidetoc","_content","Wy_wietlanieDanych","classes","affix","viewport","title","generator"],"api/WyświetlanieDanych.Program.html":["wrapper","autocollapse","logo","navbar","search","search-query","breadcrumb","sidetoggle","sidetoc","_content","Wy_wietlanieDanych_Program","Wy_wietlanieDanych_Program_syntax","methods","Wy_wietlanieDanych_Program_Main_","Wy_wietlanieDanych_Program_Main","affix","viewport","title","generator"],"toc.html":["sidetoggle","toc_filter_clear","toc_filter_input","toc","articles/toc.html","api/toc.html"],"api/toc.html":["sidetoggle","toc_filter_clear","toc_filter_input","toc",""],"articles/toc.html":["sidetoggle","toc_filter_clear","toc_filter_input","toc",""]}   P  _fileMappingG  �  {"api/WyświetlanieDanych.Form1.html":"obj/api/WyświetlanieDanych.Form1.yml","api/WyświetlanieDanych.Form2.html":"obj/api/WyświetlanieDanych.Form2.yml","api/WyświetlanieDanych.KomponentOdbieranie.html":"obj/api/WyświetlanieDanych.KomponentOdbieranie.yml","api/WyświetlanieDanych.OdbieranieDanych.html":"obj/api/WyświetlanieDanych.OdbieranieDanych.yml","api/WyświetlanieDanych.KomponentOdbieranie.Run_odbieranie.html":"obj/api/WyświetlanieDanych.KomponentOdbieranie.Run_odbieranie.yml","articles/intro.html":"articles/intro.md","index.html":"index.md","api/index.html":"api/index.md","api/WyświetlanieDanych.html":"obj/api/WyświetlanieDanych.yml","api/WyświetlanieDanych.Program.html":"obj/api/WyświetlanieDanych.Program.yml","toc.html":"toc.yml","api/toc.html":"obj/api/toc.yml","articles/toc.html":"articles/toc.md"}